`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin

        // $readmemh("sort_machine_code.mem", rom);

        for (int i = 0; i < 64; i = i + 1) begin
            rom[i] = 32'hffff_ffff;
        end

        // R-type : funct7 + rs2 + rs1 + funct3 + rd + opcode                        
        // sll -> shift left logical(논리 왼쪽 시프트) : zero extension
        // srl -> shift right logical(논리 오른쪽 시프트) : zero extension
        // sra -> shift right arithmetic(산술 오른쪽 시프트) : sign extension
        // R-type : funct7 + rs2 + rs1 + funct3 + rd + opcode      [rd] [rs1] [rs2]
        rom [0] = 32'b0000000_00100_00011_000_00000_0110011; // add  x0, x3, x4
        rom [1] = 32'b0100000_00011_00111_000_00001_0110011; // sub  x1, x7, x3
        rom [2] = 32'b0000000_00010_00100_001_00010_0110011; // sll  x2, x4, x3
        rom [3] = 32'b0000000_00011_01000_101_00011_0110011; // srl  x3, x8, x3
        rom [4] = 32'b0100000_00011_01000_101_00100_0110011; // sra  x4, x8, x3
        rom [5] = 32'b0000000_00100_00011_010_00101_0110011; // slt  x5, x3, x4
        rom [6] = 32'b0000000_00111_01000_011_00110_0110011; // sltu x6, x8, x7
        rom [7] = 32'b0000000_00100_00011_100_00111_0110011; // xor  x7, x3, x4
        rom [8] = 32'b0000000_00111_01000_110_01000_0110011; // or   x8, x8, x7
        rom [9] = 32'b0000000_00111_00100_111_01001_0110011; // and  x9, x4, x7

        //////////////////////////////////////////////////////////////////////////////////////////

        // B-type
        // beq : if(rs1 == rs2)  PC += imm
        // bne : if(rs1 != rs2)  PC += imm
        // blt : if(rs1 < rs2)   PC += imm
        // bge : if(rs1 >= rs2)  PC += imm
        // bltu : if(rs1 < rs2)  PC += imm
        // bgeu : if(rs1 >= rs2) PC += imm
        // imm[12,10:5](7bit) + rs2(5bit) + rs1(5bit) + funct3(3bit) + imm[4:1,11](5bit) + opcode(7bit)						
        // [rs1] [rs2] [imm]  
        // rom [0]  = 32'b0000000_00011_00011_000_10000_1100011; // 32'h0031_8863 - beq x3, x3, 16 (o)
        // rom [4]  = 32'b0000000_00101_00100_001_10000_1100011; // 32'h0041_9863 - bne x4, x5, 16 (o)
        // rom [8]  = 32'b1111111_11010_00010_000_00101_0010011; // 32'hffa1_8293 - addi x5, x2, -6
        // rom [12] = 32'b0000000_01000_00101_100_10000_1100011; // 32'h0082_c863 - blt x5, x8, 16 (o)
        // rom [16] = 32'b0000000_00101_00000_101_10000_1100011; // 32'h0050_5863 - bge x0, x5, 16 (o)
        // rom [20] = 32'b0000000_01010_00101_110_10000_1100011; // 32'h00a2_e863 - bltu x5, x10, 16 (x) 
        // rom [22] = 32'b0000000_00101_01000_111_10000_1100011; // 32'h0054_7863 - bgeu x8, x5, 16 (x)

        //////////////////////////////////////////////////////////////////////////////////////////

        // // S-type : imm(7bit) + rs2(5bit) + rs1(5bit) + funct3(3bit) + imm(5bit) + opcode
        // rom [0] = 32'b0000000_00011_00010_000_00010_0100011; // sb x3, 2(x2), imm = 2 , 2 + 2 = 4
        // rom [1] = 32'b0000000_00100_00010_001_01000_0100011; // sh x4, 8(x2), imm = 8 , 2 + 8 = 10
        // rom [2] = 32'b0000000_00101_00010_010_00100_0100011; // sw x5, 4(x2)  imm = 2 , 2 + 4 = 6
        // rom[0] = 32'b0000000_00101_01010_000_00000_0100011; // sb x5, 0(x10)  → data_mem[0]
        // rom[1] = 32'b0000000_00101_01010_001_00100_0100011; // sh x5, 4(x10)  → data_mem[1]
        // rom[2] = 32'b0000000_00101_01010_010_01000_0100011; // sw x5, 8(x10)  → data_mem[2]

        //////////////////////////////////////////////////////////////////////////////////////////

        // Load instructions (I-type): imm(12bit) + rs1(5bit) + funct3(3bit) + rd(5bit) + opcode(7bit)
        // IL-type
        // rom[1] = 32'b000000000000_01010_000_00010_0000011;  // lb x2, 0(x10)
        // rom[2] = 32'b000000000100_01010_001_00011_0000011;  // lh x3, 4(x10)
        // rom[3] = 32'b000000001000_01010_010_00100_0000011;  // lw x4, 8(x10)
        // rom[4] = 32'b000000000000_01010_100_00101_0000011;  // lbu x5, 0(x10)
        // rom[5] = 32'b000000000100_01010_101_00110_0000011;  // lhu x6, 4(x10)

        // I-type : imm(12bit) + rs1(5bit) + funct3(3bit) + rd(5bit) + opcode(7bit)     
        // rom[0] = 32'b000000000010_00001_000_00010_0010011; // addi x2, x1, 2      rd = rs + imm
        // rom[1] = 32'b000000000111_00001_100_00010_0010011;  // xori x2, x1, 7
        // rom[2] = 32'b000000000111_00001_110_00010_0010011;  // ori  x2, x1, 7
        // rom[3] = 32'b000000000111_00001_111_00010_0010011;  // andi x2, x1, 7
        // rom[4] = 32'b000000000011_00001_001_00010_0010011; // slli x2, x1, 3 = 8
        // rom[5] = 32'b000000000010_01000_101_00010_0010011; // srli x2, x8, 2 = 2
        // rom[6] = 32'b010000000001_01000_101_00010_0010011; // srai x2, x8, 1 = 4
        // rom[7] = 32'b000000000000_00001_010_00010_0010011; // slti x2, x1, 0  rd = (rs < imm) ? 1 : 0
        // rom[8] = 32'b111111111110_00001_011_00010_0010011; // sltiu x2, x1, -2    rd = (rs1 < imm) ? 1 : 0 (0-ex)

        //////////////////////////////////////////////////////////////////////////////////////////

        //U-Type
        //32'b imm(20bit) + rd(5bit) + opcode(7bit)
        // rom [1] = 32'b00000000000000000011_00001_0110111; // LUI x1, 3
        // rom [2] = 32'b00000000000000000011_00001_0010111; // AUIPC x1, 3

        //////////////////////////////////////////////////////////////////////////////////////////

        //J-Type
        //imm(20bit)+ rd(5bit) + opcode(7bit) c
        // imm(20bit) - imm[20,10:1,11,19:12] -> 하드웨어 단순화
        // rom[1] = 32'b0_0000001000_0_00000000_00001_1101111;  // 32'h0100_00ef - jal x1, 16 

        // //JALR(I-Type임 사실, 다음 주소 값을 레지스터에 저장 점프시킴) PC = RS1 + imm
        // //32'b imm(12bit) + rs1(5bit) + funct3(3bit) + rd(5bit) + opcode(7bit)
        // rom[15] = 32'b000000011110_00111_000_00101_1100111;  // 32'h01e3_82e7 - jalr x5, 30(x7)
    end

    assign data = rom[addr[31:2]];

endmodule

